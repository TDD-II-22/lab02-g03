`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 20.08.2022 18:46:29
// Design Name: 
// Module Name: module_key_encoding
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module module_key_encoding(
    input     logic     s1_in,
    input     logic     s0_in,
    input     logic     e1_in,
    input     logic     e2_in,
    output    logic     l0_o,
    output    logic     l1_o,
    output    logic     l2_o,
    output    logic     l3_o
    );
    
    
    
    
    
    
endmodule
